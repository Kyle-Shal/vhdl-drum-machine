library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity drum_machine is

----------WM8731 pins-----
port(AUD_BCLK: out std_logic;
AUD_XCK: out std_logic;
AUD_ADCLRCK:  out std_logic;
AUD_ADCDAT: in std_logic;
AUD_DACLRCK: out std_logic;
AUD_DACDAT: out std_logic;
---------FPGA pins-----
clock_50: in std_logic;
key: in std_logic_vector(3 downto 0);
ledr: out std_logic_vector(9 downto 0);
sw: in std_logic_vector(9 downto 0);
HEX0, HEX1, HEX2, HEX3, HEX4, HEX5 : out std_logic_vector (6 downto 0);
FPGA_I2C_SCLK: out std_logic;
FPGA_I2C_SDAT: inout std_logic );

end drum_machine;


architecture logic of drum_machine is

signal aud_mono: std_logic_vector(31 downto 0):=(others=>'0');
signal read_addr: integer range 0 to 256000:=0;
signal ROM_ADDR: std_logic_vector(17 downto 0);
signal ROM_OUT: std_logic_vector(15 downto 0);
signal clock_12pll: std_logic;
signal config_busy: std_logic;
signal config_done: std_logic;
signal config_send_flag: std_logic;
signal config_data: std_logic_vector(15 downto 0);
signal DA_CLR: std_logic:='0';
signal k0_sig, k1_sig, k2_sig, k3_sig: std_logic := '0';
signal DISP0, DISP1, DISP2, DISP3, DISP4, DISP5: std_logic_vector (4 downto 0) := "11111";
signal config_count: integer range 0 to 7:=0;
    
	 component pll is
        port (
            clk_clk                         : in  std_logic                     := 'X';             -- clk
            clock_12_clk                    : out std_logic;                                        -- clk
            reset_reset_n                   : in  std_logic                     := 'X';             -- reset_n
            onchip_memory2_0_s1_address     : in  std_logic_vector(17 downto 0) := (others => 'X'); -- address
            onchip_memory2_0_s1_debugaccess : in  std_logic                     := 'X';             -- debugaccess
            onchip_memory2_0_s1_clken       : in  std_logic                     := 'X';             -- clken
            onchip_memory2_0_s1_chipselect  : in  std_logic                     := 'X';             -- chipselect
            onchip_memory2_0_s1_write       : in  std_logic                     := 'X';             -- write
            onchip_memory2_0_s1_readdata    : out std_logic_vector(15 downto 0);                    -- readdata
            onchip_memory2_0_s1_writedata   : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
            onchip_memory2_0_s1_byteenable  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
		      onchip_memory2_0_reset1_reset   : in  std_logic                     := 'X'              -- reset		
        );
		  end component pll;

component audio_data is
	port (clock_12: in std_logic;
		bclk: out std_logic;
		daclr: out std_logic;
		dacdat: out std_logic;
		data_in: in std_logic_vector(31 downto 0));
end component audio_data;





component audio_config is
	port( busy_flag: out std_logic;
		sclk: out std_logic;
		send_flag: in std_logic;
		sdin: inout std_logic;
		done_flag: out std_logic;
		data_in: in std_logic_vector(15 downto 0);
		clock_50_in: in std_logic );
end component audio_config;
 
 component seven_segment_decoder is
	port(input: in std_logic_vector(4 downto 0);
		  output: out std_logic_vector(6 downto 0));
 end component;
 

begin

--- on chip memory component generated by Qsys
 u0 : component pll
        port map (
            clk_clk       => clock_50,                                           -- clk.clk
            reset_reset_n => '1',                                                -- reset.reset_n
            clock_12_clk  => clock_12pll, 												   -- clock_12.clk
				onchip_memory2_0_s1_address     => ROM_ADDR,
            onchip_memory2_0_s1_debugaccess =>'0',                               -- debugaccess
            onchip_memory2_0_s1_clken       =>'1',                               -- clken
            onchip_memory2_0_s1_chipselect  =>'1',                               -- chipselect
            onchip_memory2_0_s1_write      =>'0',                                -- write
            onchip_memory2_0_s1_readdata   =>ROM_OUT,                            -- readdata
            onchip_memory2_0_s1_writedata  =>(others=>'0'),
            onchip_memory2_0_s1_byteenable  =>"11",
				onchip_memory2_0_reset1_reset=>'0'
				);
				

audio_data_sender: component audio_data port map(clock_12pll, AUD_BCLK, DA_CLR, AUD_DACDAT, aud_mono);
audio_configuration: component audio_config port map(config_busy, FPGA_I2C_SCLK, config_send_flag, FPGA_I2C_SDAT, config_done, config_data, clock_50);

HEXDISP0: component seven_segment_decoder port map (DISP0,HEX0);
HEXDISP1: component seven_segment_decoder port map (DISP1,HEX1);
HEXDISP2: component seven_segment_decoder port map (DISP2,HEX2);
HEXDISP3: component seven_segment_decoder port map (DISP3,HEX3);
HEXDISP4: component seven_segment_decoder port map (DISP4,HEX4);
HEXDISP5: component seven_segment_decoder port map (DISP5,HEX5);

AUD_XCK<=clock_12pll;
AUD_DACLRCK<=DA_CLR;
	
ROM_ADDR<=std_logic_vector(to_unsigned(read_addr,18));

process (clock_12pll)
begin

if rising_edge(clock_12pll)then

 	if(SW(9)='0' or (k0_sig = '0' and k1_sig = '0' and k2_sig = '0' and k3_sig = '0'))then --- Idle State
	read_addr<=0;
	aud_mono<=(others=>'0');
	else --- Output audio
	aud_mono(15 downto 0)<=ROM_OUT;
	aud_mono(31 downto 16)<=ROM_OUT;
	  if(DA_CLR='1' and k0_sig = '1')then
			if(read_addr<28325)then
				read_addr<=read_addr+1;
			else
				read_addr<=0;
				k0_sig<='0';
			end if;
		elsif(DA_CLR='1' and k1_sig = '1')then
			if(read_addr<44416)then
				read_addr<=read_addr+1;
			else
				read_addr<=0;
				k1_sig<='0';
			end if;
		elsif(DA_CLR='1' and k2_sig = '1')then
			if(read_addr<58878)then
				read_addr<=read_addr+1;
			else
				read_addr<=0;
				k2_sig<='0';
			end if;
		elsif(DA_CLR='1' and k3_sig = '1')then
			if(read_addr<68863)then
				read_addr<=read_addr+1;
			else
				read_addr<=0;
				k3_sig<='0';
			end if;
		end if;
	end if;

	if (KEY(0)='0' AND SW(9)='1') then --- Hi Hat
		read_addr<=0;
		aud_mono<=(others=>'0');
		k0_sig <= '1';
		k1_sig <= '0';
		k2_sig <= '0';
		k3_sig <= '0';
  		DISP5 <= "01010"; ---H
		DISP4 <= "01011"; ---I
		DISP3 <= "11111"; ---
		DISP2 <= "01010"; ---H
		DISP1 <= "00101"; ---A
		DISP0 <= "10001"; ---t
		
	elsif(KEY(1)='0' AND SW(9)='1') then --- Percussion
		read_addr<=28326;
		aud_mono<=(others=>'0');
		k0_sig <= '0';
		k1_sig <= '1';
		k2_sig <= '0';
		k3_sig <= '0';
		DISP5 <= "01110"; ---P
		DISP4 <= "01001"; ---E
		DISP3 <= "01111"; ---r
		DISP2 <= "00111"; ---c
		DISP1 <= "11111"; ---
		DISP0 <= "11111"; ---
		
	elsif(KEY(2)='0' AND SW(9)='1') then --- Bass
		read_addr<=44417;
		aud_mono<=(others=>'0');
		k0_sig <= '0';
		k1_sig <= '0';
		k2_sig <= '1';
		k3_sig <= '0';
		DISP5 <= "00110"; ---b
		DISP4 <= "00101"; ---A
		DISP3 <= "10000"; ---S
		DISP2 <= "10000"; ---S
		DISP1 <= "11111"; ---
		DISP0 <= "11111"; ---
		
	elsif(KEY(3)='0' AND SW(9)='1') then --- Snare
		read_addr<=58879;
		aud_mono<=(others=>'0');
		k0_sig <= '0';
		k1_sig <= '0';
		k2_sig <= '0';
		k3_sig <= '1';
		DISP5 <= "10000"; ---S
		DISP4 <= "01101"; ---n
		DISP3 <= "00101"; ---A
		DISP2 <= "01111"; ---r
		DISP1 <= "01001"; ---E
		DISP0 <= "11111"; ---
	elsif(SW(9)='1') then
		DISP5 <= "01000"; ---d
		DISP4 <= "01111"; ---r
		DISP3 <= "10010"; ---u
		DISP2 <= "01100"; ---M
		DISP1 <= "10000"; ---S
		DISP0 <= "11111"; ---
		LEDR(config_count) <= '1';
	end if;
	
	if(SW(9)='0' and KEY(0)='0') then
		DISP5 <= "10011"; ---V
		DISP4 <= "00000"; ---O
		DISP3 <= "10100"; ---L
		DISP2 <= "00001"; ---1
		DISP1 <= "11111"; ---
		DISP0 <= "11111"; ---
	elsif(SW(9)='0' and KEY(1)='0') then
		DISP5 <= "10011"; ---V
		DISP4 <= "00000"; ---O
		DISP3 <= "10100"; ---L
		DISP2 <= "00010"; ---2
		DISP1 <= "11111"; ---
		DISP0 <= "11111"; ---
	elsif(SW(9)='0' and KEY(2)='0') then
		DISP5 <= "10011"; ---V
		DISP4 <= "00000"; ---O
		DISP3 <= "10100"; ---L
		DISP2 <= "00011"; ---3
		DISP1 <= "11111"; ---
		DISP0 <= "11111"; ---
	elsif(SW(9)='0' and KEY(3)='0') then
		DISP5 <= "10011"; ---V
		DISP4 <= "00000"; ---O
		DISP3 <= "10100"; ---L
		DISP2 <= "00100"; ---4
		DISP1 <= "11111"; ---
		DISP0 <= "11111"; ---
	elsif(SW(9)='0') then
		DISP5 <= "10011"; ---V
		DISP4 <= "00000"; ---O
		DISP3 <= "10100"; ---L
		DISP2 <= "10010"; ---u
		DISP1 <= "01100"; ---M
		DISP0 <= "01001"; ---E
	end if;
end if;

end process;	

process (clock_50)
begin

 if rising_edge(clock_50) then
		
		config_send_flag<='0';
		
		if config_busy='0' then
			if (SW(9)='0' AND KEY(0)='0') then --- VOL1 (-15dB)
			config_data(15 downto 9)<="0000010";
			config_data(8 downto 0)<="101101010";
			config_send_flag<='1';
			
			elsif (SW(9)='0' AND KEY(1)='0') then --- VOL2 (-8dB)
			config_data(15 downto 9)<="0000010";
			config_data(8 downto 0)<="101110001";
			config_send_flag<='1';
			
			elsif (SW(9)='0' AND KEY(2)='0') then --- VOL3 (-1dB)
			config_data(15 downto 9)<="0000010";
			config_data(8 downto 0)<="101111000";
			config_send_flag<='1';
		
			elsif (SW(9)='0' AND KEY(3)='0') then --- VOL4 (+6dB)
			config_data(15 downto 9)<="0000010";
			config_data(8 downto 0)<="101111111";
			config_send_flag<='1';
			
			elsif ((config_count=0 and config_done = '1') or (SW(0)='1' and SW(1) = '0')) then --- Activate control interface
			config_data(15 downto 9)<="0001001";
			config_data(8 downto 0)<="111111111";
			config_send_flag<='1';
			config_count <= config_count + 1 ;
			
			elsif ((config_count=1 and config_done = '1') or (SW(0)='0' and SW(1) = '1')) then --- Turn off Line Input, Microphone Input, and ADC to conserve power
			config_data(15 downto 9)<="0000110";
			config_data(8 downto 0)<="000000111";
			config_send_flag<='1';
			config_count <= config_count + 1 ;		
			
			elsif ((config_count=2 and config_done = '1') or (SW(0)='1' and SW(1) = '1')) then --- Set DSP/PCM mode with MSB available on 2nd BCLK rising edge, 16 bit mode, and slave mode
			config_data(15 downto 9)<="0000111"; 
			config_data(8 downto 0)<="000010011";	
			config_send_flag<='1';
			config_count <= config_count + 1 ;	
			
			elsif ((config_count=3 and config_done = '1') or (SW(2)='1' and SW(3) = '0')) then --- Set USB mode 250 fs base oversampling rate
			config_data(15 downto 9)<="0001000";
			config_data(8 downto 0)<="000000001";
			config_send_flag<='1';
			config_count <= config_count + 1 ;		
				
			elsif ((config_count=4 and config_done = '1') or (SW(2)='0' and SW(3) = '1')) then --- Enable DAC to LINOUT and Disable Mic
			config_data(15 downto 9)<="0000100";
			config_data(8 downto 0)<="000010010";
			config_send_flag<='1';
			config_count <= config_count + 1 ;		
			
			elsif ((config_count=5 and config_done = '1') or (SW(2)='1' and SW(3) = '1')) then --- Disable DAC soft mute
			config_data(15 downto 9)<="0000101";
			config_data(8 downto 0)<="000000000";
			config_send_flag<='1';
			config_count <= config_count + 1 ;		
			
			elsif((config_count=6 and config_done = '1')) then --- Set Volume to level 4 (+6dB)
			config_data(15 downto 9)<="0000010";
			config_data(8 downto 0)<="101111111";
			config_send_flag<='1';
			config_count <= config_count + 1 ;		
			end if;
		end if;
 end if;
end process;
end logic;